----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:02:11 07/18/2023 
-- Design Name: 
-- Module Name:    decode_select_ins - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity decode_select_ins is
	port(
		i: in  STD_LOGIC_VECTOR(1 downto 0);
		o: out STD_LOGIC_VECTOR(3 downto 0));
end decode_select_ins;

architecture Behavioral of decode_select_ins is
begin
	with i select
	o <= 	"0001" when "00",
			"0010" when "01",
			"0100" when "10",
			"1000" when others;
			

end Behavioral;

